//////////////////////////////////////////////////////////////////
///
/// Project Name: 	avalon_enforcer
///
/// File Name: 		general_pack.sv
///
//////////////////////////////////////////////////////////////////
///
/// Author: 		Ariel Kalish
///
/// Date Created: 	19.3.2020
///
/// Company: 		----
///
//////////////////////////////////////////////////////////////////
///
/// Description: 	Package containing general functions
///
//////////////////////////////////////////////////////////////////

package general_pack;

	function int log2up_func (int num);
		if (num == 1) begin
			return 1;
		end else begin
			return $clog2(num);
		end
	endfunction

endpackage

